module UART_Handshake();
endmodule